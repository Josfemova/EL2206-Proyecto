* NGSPICE file created from nand_Lpnx2.ext - technology: scmos

.option scale=0.09u

M1000 vdd in out vdd pfet w=8 l=4
+  ad=48 pd=28 as=80 ps=52
M1001 out in a_n1_n9# Gnd nfet w=4 l=4
+  ad=20 pd=18 as=24 ps=20
M1002 a_n1_n9# in Gnd Gnd nfet w=4 l=4
+  ad=0 pd=0 as=20 ps=18
M1003 out in vdd vdd pfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
C0 Gnd in 0.04fF
C1 out Gnd 0.08fF
C2 out in 0.23fF
C3 vdd in 0.45fF
C4 out vdd 0.52fF
C5 Gnd 0 0.10fF $ **FLOATING
C6 out 0 0.26fF $ **FLOATING
C7 in 0 0.44fF $ **FLOATING
C8 vdd 0 0.61fF $ **FLOATING
