* NGSPICE file created from nand_Wpnx3.ext - technology: scmos

.option scale=0.09u

M1000 out in a_n1_n17# Gnd nfet w=12 l=2
+  ad=60 pd=34 as=72 ps=36
M1001 vdd in out vdd pfet w=24 l=2
+  ad=144 pd=60 as=240 ps=116
M1002 out in vdd vdd pfet w=24 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_n1_n17# in Gnd Gnd nfet w=12 l=2
+  ad=0 pd=0 as=60 ps=34
C0 in vdd 0.32fF
C1 Gnd in 0.03fF
C2 out vdd 1.02fF
C3 Gnd out 0.08fF
C4 in out 0.11fF
C5 Gnd 0 0.11fF $ **FLOATING
C6 out 0 0.31fF $ **FLOATING
C7 in 0 0.37fF $ **FLOATING
C8 vdd 0 0.91fF $ **FLOATING
