* NGSPICE file created from nand_Lnx3.ext - technology: scmos

.option scale=0.09u

M1000 vdd in out vdd pfet w=8 l=2
+  ad=48 pd=28 as=128 ps=100
M1001 a_0_n9# in out Gnd nfet w=4 l=6
+  ad=16 pd=16 as=20 ps=18
M1002 a_10_n9# in a_0_n9# Gnd nfet w=4 l=6
+  ad=20 pd=18 as=0 ps=0
M1003 out in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd in 0.33fF
C1 vdd out 0.57fF
C2 in out 0.06fF
C3 a_10_n9# out 0.08fF
C4 a_10_n9# 0 0.01fF $ **FLOATING
C5 out 0 0.38fF $ **FLOATING
C6 in 0 0.47fF $ **FLOATING
C7 vdd 0 0.64fF $ **FLOATING
