* NGSPICE file created from nand_Wpnx2.ext - technology: scmos

.option scale=0.09u

M1000 vdd in out vdd pfet w=16 l=2
+  ad=96 pd=44 as=160 ps=84
M1001 a_n1_n13# in Gnd Gnd nfet w=8 l=2
+  ad=48 pd=28 as=40 ps=26
M1002 out in a_n1_n13# Gnd nfet w=8 l=2
+  ad=40 pd=26 as=0 ps=0
M1003 out in vdd vdd pfet w=16 l=2
+  ad=0 pd=0 as=0 ps=0
C0 Gnd out 0.08fF
C1 vdd in 0.33fF
C2 Gnd in 0.03fF
C3 vdd out 0.81fF
C4 in out 0.11fF
C5 Gnd 0 0.11fF $ **FLOATING
C6 out 0 0.28fF $ **FLOATING
C7 in 0 0.37fF $ **FLOATING
C8 vdd 0 0.72fF $ **FLOATING
