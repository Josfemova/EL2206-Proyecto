* NGSPICE file created from nand_Lnx3.ext - technology: scmos

.option scale=0.09u

M1000 vdd in out vdd pfet w=8 l=2
+  ad=48 pd=28 as=80 ps=52
M1001 a_0_n9# in Gnd Gnd nfet w=4 l=6
+  ad=16 pd=16 as=20 ps=18
M1002 out in a_0_n9# Gnd nfet w=4 l=6
+  ad=20 pd=18 as=0 ps=0
M1003 out in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in out 0.03fF
C1 Gnd in 0.03fF
C2 vdd in 0.33fF
C3 Gnd out 0.05fF
C4 vdd out 0.56fF
C5 Gnd 0 0.13fF $ **FLOATING
C6 out 0 0.26fF $ **FLOATING
C7 in 0 0.47fF $ **FLOATING
C8 vdd 0 0.64fF $ **FLOATING
