magic
tech scmos
timestamp 1667800846
<< nwell >>
rect -14 1 21 26
<< ntransistor >>
rect -3 -33 -1 -29
rect 5 -33 7 -29
<< ptransistor >>
rect -3 7 -1 15
rect 5 7 7 15
<< ndiffusion >>
rect -4 -33 -3 -29
rect -1 -33 5 -29
rect 7 -33 8 -29
<< pdiffusion >>
rect -4 7 -3 15
rect -1 7 0 15
rect 4 7 5 15
rect 7 7 8 15
<< ndcontact >>
rect -8 -33 -4 -29
rect 8 -33 12 -29
<< pdcontact >>
rect -8 7 -4 15
rect 0 7 4 15
rect 8 7 12 15
<< psubstratepcontact >>
rect -8 -41 -4 -37
rect 0 -41 4 -37
rect 8 -41 12 -37
<< nsubstratencontact >>
rect -8 19 -4 23
rect 0 19 4 23
rect 8 19 12 23
<< polysilicon >>
rect -3 15 -1 27
rect 5 15 7 27
rect -3 -29 -1 7
rect 5 -29 7 7
rect 15 -9 17 27
rect -3 -43 -1 -33
rect 5 -43 7 -33
rect 15 -43 17 -13
<< polycontact >>
rect -4 27 0 31
rect 4 27 8 31
rect 14 27 18 31
rect 14 -13 18 -9
<< metal1 >>
rect -4 31 8 35
rect 14 31 18 35
rect -14 19 -8 23
rect -4 19 0 23
rect 4 19 8 23
rect 12 19 21 23
rect 0 15 4 19
rect -8 -9 -4 7
rect 8 -9 12 7
rect -8 -13 14 -9
rect -8 -37 -4 -33
rect -14 -41 -8 -37
rect -4 -41 0 -37
rect 4 -41 8 -37
rect 12 -41 21 -37
<< labels >>
rlabel metal1 14 31 18 35 6 out
rlabel metal1 0 31 4 35 5 in
rlabel metal1 -14 19 -10 23 3 vdd
rlabel metal1 -14 -41 -10 -37 2 Gnd
<< end >>
