* NGSPICE file created from nand_distcompx2.ext - technology: scmos

.option scale=0.09u

M1000 out in vdd vdd pfet w=8 l=2
+  ad=80 pd=52 as=96 ps=40
M1001 vdd in out vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 out in a_n4_n9# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=48 ps=32
M1003 a_n4_n9# in Gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
C0 in Gnd 0.03fF
C1 Gnd out 0.08fF
C2 in vdd 0.37fF
C3 vdd out 0.69fF
C4 in out 0.11fF
C5 Gnd 0 0.13fF $ **FLOATING
C6 out 0 0.27fF $ **FLOATING
C7 in 0 0.39fF $ **FLOATING
C8 vdd 0 0.65fF $ **FLOATING
