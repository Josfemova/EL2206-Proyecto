magic
tech scmos
timestamp 1667810131
<< nwell >>
rect -20 1 27 26
<< ntransistor >>
rect -9 -9 -7 -5
rect 11 -9 13 -5
<< ptransistor >>
rect -9 7 -7 15
rect 11 7 13 15
<< ndiffusion >>
rect -10 -9 -9 -5
rect -7 -9 11 -5
rect 13 -9 14 -5
<< pdiffusion >>
rect -10 7 -9 15
rect -7 7 -6 15
rect 10 7 11 15
rect 13 7 14 15
<< ndcontact >>
rect -14 -9 -10 -5
rect 14 -9 18 -5
<< pdcontact >>
rect -14 7 -10 15
rect -6 7 10 15
rect 14 7 18 15
<< psubstratepcontact >>
rect -16 -17 -12 -13
rect -4 -17 0 -13
rect 4 -17 8 -13
rect 15 -17 19 -13
<< nsubstratencontact >>
rect -17 19 -13 23
rect -4 19 0 23
rect 4 19 8 23
rect 15 19 19 23
<< polysilicon >>
rect -9 15 -7 27
rect 11 15 13 27
rect -9 -5 -7 7
rect 11 -5 13 7
rect 21 3 23 27
rect -9 -19 -7 -9
rect 11 -19 13 -9
rect 21 -19 23 -1
<< polycontact >>
rect -10 27 -6 31
rect 10 27 14 31
rect 20 27 24 31
rect 20 -1 24 3
<< metal1 >>
rect -10 31 14 35
rect 20 31 24 35
rect -20 19 -17 23
rect -13 19 -4 23
rect 0 15 4 23
rect 8 19 15 23
rect 19 19 27 23
rect -14 3 -10 7
rect 14 3 18 7
rect -14 -1 20 3
rect 14 -5 18 -1
rect -14 -13 -10 -9
rect -20 -17 -16 -13
rect -12 -17 -4 -13
rect 0 -17 4 -13
rect 8 -17 15 -13
rect 19 -17 24 -13
<< labels >>
rlabel metal1 -17 -17 -13 -13 2 Gnd
rlabel metal1 -17 19 -13 23 3 vdd
rlabel metal1 20 31 24 35 6 out
rlabel metal1 0 31 4 35 5 in
<< end >>
