Sim file

.INCLUDE "tsmc018.lib"
.INCLUDE "nand_Wnx3.spice"

V1 vdd Gnd 1.8
V2 in Gnd PULSE(0 1.8 0.05n 0.1f 0.1f 0.6n 1.2n)

.MEAS TRAN tphl TRIG V(in) VAL=0.9 RISE=1 
+               TARG V(out) VAL=0.9 FALL=1
.MEAS TRAN tplh TRIG V(in) VAL=0.9 FALL=1 
+               TARG V(out) VAL=0.9 RISE=1


.MEAS TRAN tpd PARAM=(tphl+tplh)/2

.MEAS TRAN corriente_max MAX I(V1)
.MEAS TRAN pmax PARAM=corriente_max*1.8

.TRAN 10p 1.2n 

.end
