magic
tech scmos
timestamp 1667804431
<< nwell >>
rect -17 1 22 26
<< ntransistor >>
rect -5 -9 -1 -5
rect 5 -9 9 -5
<< ptransistor >>
rect -5 7 -1 15
rect 5 7 9 15
<< ndiffusion >>
rect -6 -9 -5 -5
rect -1 -9 5 -5
rect 9 -9 10 -5
<< pdiffusion >>
rect -6 7 -5 15
rect -1 7 0 15
rect 4 7 5 15
rect 9 7 10 15
<< ndcontact >>
rect -10 -9 -6 -5
rect 10 -9 14 -5
<< pdcontact >>
rect -10 7 -6 15
rect 0 7 4 15
rect 10 7 14 15
<< psubstratepcontact >>
rect -10 -17 -6 -13
rect 0 -17 4 -13
rect 10 -17 14 -13
<< nsubstratencontact >>
rect -10 19 -6 23
rect 0 19 4 23
rect 10 19 14 23
<< polysilicon >>
rect -5 15 -1 27
rect 5 15 9 27
rect -5 -5 -1 7
rect 5 -5 9 7
rect 16 3 18 27
rect -5 -19 -1 -9
rect 5 -19 9 -9
rect 16 -19 18 -1
<< polycontact >>
rect -5 27 -1 31
rect 5 27 9 31
rect 15 27 19 31
rect 15 -1 19 3
<< metal1 >>
rect -5 31 9 35
rect 15 31 19 35
rect -17 19 -10 23
rect -6 19 0 23
rect 4 19 10 23
rect 14 19 22 23
rect 0 15 4 19
rect -10 3 -6 7
rect 10 3 14 7
rect -10 -1 15 3
rect 10 -5 14 -1
rect -10 -13 -6 -9
rect -17 -17 -10 -13
rect -6 -17 0 -13
rect 4 -17 10 -13
rect 14 -17 20 -13
<< labels >>
rlabel metal1 0 31 4 35 5 in
rlabel metal1 -14 19 -10 23 3 vdd
rlabel metal1 -15 -17 -11 -13 2 Gnd
rlabel metal1 15 31 19 35 6 out
<< end >>
