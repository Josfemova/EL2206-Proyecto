* NGSPICE file created from nand_dist_nmos-pmosx3.ext - technology: scmos

.option scale=0.09u

M1000 a_n1_n33# in Gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1001 a_7_n33# in a_n1_n33# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1002 vdd in out vdd pfet w=8 l=2
+  ad=48 pd=28 as=80 ps=52
M1003 out in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in vdd 0.33fF
C1 out vdd 0.49fF
C2 Gnd in 0.03fF
C3 a_7_n33# Gnd 0.02fF
C4 out Gnd 0.01fF
C5 out in 0.11fF
C6 a_7_n33# 0 0.01fF $ **FLOATING
C7 Gnd 0 0.11fF $ **FLOATING
C8 out 0 0.48fF $ **FLOATING
C9 in 0 0.65fF $ **FLOATING
C10 vdd 0 0.55fF $ **FLOATING
