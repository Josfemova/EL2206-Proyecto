magic
tech scmos
timestamp 1667799124
<< nwell >>
rect -14 1 21 26
<< ntransistor >>
rect -3 -9 -1 -5
rect 5 -9 7 -5
<< ptransistor >>
rect -3 7 -1 15
rect 5 7 7 15
<< ndiffusion >>
rect -4 -9 -3 -5
rect -1 -9 5 -5
rect 7 -9 8 -5
<< pdiffusion >>
rect -4 7 -3 15
rect -1 7 0 15
rect 4 7 5 15
rect 7 7 8 15
<< ndcontact >>
rect -8 -9 -4 -5
rect 8 -9 12 -5
<< pdcontact >>
rect -8 7 -4 15
rect 0 7 4 15
rect 8 7 12 15
<< psubstratepcontact >>
rect -8 -17 -4 -13
rect 0 -17 4 -13
rect 8 -17 12 -13
<< nsubstratencontact >>
rect -8 19 -4 23
rect 0 19 4 23
rect 8 19 12 23
<< polysilicon >>
rect -3 15 -1 27
rect 5 15 7 27
rect -3 -5 -1 7
rect 5 -5 7 7
rect 15 3 17 27
rect -3 -19 -1 -9
rect 5 -19 7 -9
rect 15 -19 17 -1
<< polycontact >>
rect -4 27 0 31
rect 4 27 8 31
rect 14 27 18 31
rect 14 -1 18 3
<< metal1 >>
rect -4 31 8 35
rect 14 31 18 35
rect -14 19 -8 23
rect -4 19 0 23
rect 4 19 8 23
rect 12 19 21 23
rect 0 15 4 19
rect -8 3 -4 7
rect 8 3 12 7
rect -8 -1 14 3
rect 8 -5 12 -1
rect -8 -13 -4 -9
rect -14 -17 -8 -13
rect -4 -17 0 -13
rect 4 -17 8 -13
rect 12 -17 21 -13
<< labels >>
rlabel metal1 -14 -17 -10 -13 2 Gnd
rlabel metal1 14 31 18 35 6 out
rlabel metal1 0 31 4 35 5 in
rlabel metal1 -14 19 -10 23 3 vdd
<< end >>
