magic
tech scmos
timestamp 1667801468
<< nwell >>
rect -14 1 21 26
<< ntransistor >>
rect -3 -13 -1 -5
rect 5 -13 7 -5
<< ptransistor >>
rect -3 7 -1 15
rect 5 7 7 15
<< ndiffusion >>
rect -4 -13 -3 -5
rect -1 -13 5 -5
rect 7 -13 8 -5
<< pdiffusion >>
rect -4 7 -3 15
rect -1 7 0 15
rect 4 7 5 15
rect 7 7 8 15
<< ndcontact >>
rect -8 -13 -4 -5
rect 8 -13 12 -5
<< pdcontact >>
rect -8 7 -4 15
rect 0 7 4 15
rect 8 7 12 15
<< psubstratepcontact >>
rect -8 -21 -4 -17
rect 0 -21 4 -17
rect 8 -21 12 -17
<< nsubstratencontact >>
rect -8 19 -4 23
rect 0 19 4 23
rect 8 19 12 23
<< polysilicon >>
rect -3 15 -1 27
rect 5 15 7 27
rect -3 -5 -1 7
rect 5 -5 7 7
rect 15 3 17 27
rect -3 -23 -1 -13
rect 5 -23 7 -13
rect 15 -23 17 -1
<< polycontact >>
rect -4 27 0 31
rect 4 27 8 31
rect 14 27 18 31
rect 14 -1 18 3
<< metal1 >>
rect -4 31 8 35
rect 14 31 18 35
rect -14 19 -8 23
rect -4 19 0 23
rect 4 19 8 23
rect 12 19 21 23
rect 0 15 4 19
rect -8 3 -4 7
rect 8 3 12 7
rect -8 -1 14 3
rect -8 -5 -4 -1
rect 8 -5 12 -1
rect -8 -17 -4 -13
rect -14 -21 -8 -17
rect -4 -21 0 -17
rect 4 -21 8 -17
rect 12 -21 21 -17
<< labels >>
rlabel metal1 14 31 18 35 6 out
rlabel metal1 0 31 4 35 5 in
rlabel metal1 -14 19 -10 23 3 vdd
rlabel metal1 -14 -21 -10 -17 2 Gnd
<< end >>
