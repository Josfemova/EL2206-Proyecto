* NGSPICE file created from nand_dist_nmos-pmosx2.ext - technology: scmos

.option scale=0.09u

M1000 vdd in Gnd vdd pfet w=8 l=2
+  ad=48 pd=28 as=128 ps=100
M1001 a_n1_n21# in Gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=40 ps=36
M1002 Gnd in a_n1_n21# Gnd nfet w=4 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Gnd in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in vdd 0.33fF
C1 Gnd vdd 0.49fF
C2 Gnd a_15_n31# 0.02fF
C3 in Gnd 0.14fF
C4 a_15_n31# 0 0.02fF
C5 Gnd 0 0.51fF $ **FLOATING
C6 in 0 0.51fF $ **FLOATING
C7 vdd 0 0.55fF $ **FLOATING
