* NGSPICE file created from nand_dist_nmos-pmosx2.ext - technology: scmos

.option scale=0.09u

M1000 vdd in out vdd pfet w=8 l=2
+  ad=48 pd=28 as=80 ps=52
M1001 a_n1_n21# in Gnd Gnd nfet w=4 l=2
+  ad=24 pd=20 as=20 ps=18
M1002 out in a_n1_n21# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1003 out in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 out in 0.11fF
C1 out vdd 0.49fF
C2 out Gnd 0.04fF
C3 in vdd 0.33fF
C4 in Gnd 0.03fF
C5 Gnd 0 0.11fF $ **FLOATING
C6 out 0 0.41fF $ **FLOATING
C7 in 0 0.51fF $ **FLOATING
C8 vdd 0 0.55fF $ **FLOATING
