magic
tech scmos
timestamp 1667804867
<< nwell >>
rect -22 1 24 26
<< ntransistor >>
rect -7 -9 -1 -5
rect 5 -9 11 -5
<< ptransistor >>
rect -7 7 -1 15
rect 5 7 11 15
<< ndiffusion >>
rect -8 -9 -7 -5
rect -1 -9 5 -5
rect 11 -9 12 -5
<< pdiffusion >>
rect -8 7 -7 15
rect -1 7 0 15
rect 4 7 5 15
rect 11 7 12 15
<< ndcontact >>
rect -12 -9 -8 -5
rect 12 -9 16 -5
<< pdcontact >>
rect -12 7 -8 15
rect 0 7 4 15
rect 12 7 16 15
<< psubstratepcontact >>
rect -12 -17 -8 -13
rect 0 -17 4 -13
rect 12 -17 16 -13
<< nsubstratencontact >>
rect -12 19 -8 23
rect 0 19 4 23
rect 13 19 17 23
<< polysilicon >>
rect -7 15 -1 27
rect 5 15 11 27
rect -7 -5 -1 7
rect 5 -5 11 7
rect 18 3 20 27
rect -7 -19 -1 -9
rect 5 -19 11 -9
rect 18 -19 20 -1
<< polycontact >>
rect -7 27 -1 31
rect 5 27 11 31
rect 17 27 21 31
rect 17 -1 21 3
<< metal1 >>
rect -7 31 11 35
rect 17 31 21 35
rect -22 19 -12 23
rect -8 19 0 23
rect 4 19 13 23
rect 17 19 24 23
rect 0 15 4 19
rect -12 3 -8 7
rect 12 3 16 7
rect -12 -1 17 3
rect -12 -2 16 -1
rect 12 -5 16 -2
rect -12 -13 -8 -9
rect -22 -17 -12 -13
rect -8 -17 0 -13
rect 4 -17 12 -13
rect 16 -17 24 -13
<< labels >>
rlabel metal1 0 31 4 35 5 in
rlabel metal1 -14 19 -10 23 3 vdd
rlabel metal1 -15 -17 -11 -13 2 Gnd
rlabel metal1 17 31 21 35 6 out
<< end >>
