magic
tech scmos
timestamp 1667803821
<< nwell >>
rect -14 1 21 43
<< ntransistor >>
rect -3 -17 -1 -5
rect 5 -17 7 -5
<< ptransistor >>
rect -3 7 -1 31
rect 5 7 7 31
<< ndiffusion >>
rect -4 -17 -3 -5
rect -1 -17 5 -5
rect 7 -17 8 -5
<< pdiffusion >>
rect -4 7 -3 31
rect -1 7 0 31
rect 4 7 5 31
rect 7 7 8 31
<< ndcontact >>
rect -8 -17 -4 -5
rect 8 -17 12 -5
<< pdcontact >>
rect -8 7 -4 31
rect 0 7 4 31
rect 8 7 12 31
<< psubstratepcontact >>
rect -8 -25 -4 -21
rect 0 -25 4 -21
rect 8 -25 12 -21
<< nsubstratencontact >>
rect -8 35 -4 39
rect 0 35 4 39
rect 8 35 12 39
<< polysilicon >>
rect -3 31 -1 44
rect 5 31 7 44
rect -3 -5 -1 7
rect 5 -5 7 7
rect 15 3 17 44
rect -3 -27 -1 -17
rect 5 -27 7 -17
rect 15 -27 17 -1
<< polycontact >>
rect -4 44 0 48
rect 4 44 8 48
rect 14 44 18 48
rect 14 -1 18 3
<< metal1 >>
rect -4 48 8 52
rect 14 48 18 52
rect -14 35 -8 39
rect -4 35 0 39
rect 4 35 8 39
rect 12 35 21 39
rect 0 31 4 35
rect -8 3 -4 7
rect 8 3 12 7
rect -8 -1 14 3
rect 8 -5 12 -1
rect -8 -21 -4 -17
rect -14 -25 -8 -21
rect -4 -25 0 -21
rect 4 -25 8 -21
rect 12 -25 21 -21
<< labels >>
rlabel metal1 -14 -25 -10 -21 2 Gnd
rlabel metal1 14 48 18 52 6 out
rlabel metal1 0 48 4 52 5 in
rlabel metal1 -14 35 -10 39 3 vdd
<< end >>
