* NGSPICE file created from nand_Wnx2.ext - technology: scmos

.option scale=0.09u

M1000 vdd in Gnd vdd pfet w=8 l=2
+  ad=48 pd=28 as=128 ps=100
M1001 a_n1_n13# in Gnd Gnd nfet w=8 l=2
+  ad=48 pd=28 as=80 ps=52
M1002 Gnd in a_n1_n13# Gnd nfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Gnd in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd Gnd 0.58fF
C1 Gnd in 0.14fF
C2 vdd in 0.33fF
C3 Gnd 0 0.40fF $ **FLOATING
C4 in 0 0.37fF $ **FLOATING
C5 vdd 0 0.55fF $ **FLOATING
