* NGSPICE file created from nand_referencia.ext - technology: scmos

.option scale=0.09u

M1000 vdd in out vdd pfet w=8 l=2
+  ad=48 pd=28 as=80 ps=52
M1001 out in a_n1_n9# Gnd nfet w=4 l=2
+  ad=20 pd=18 as=24 ps=20
M1002 a_n1_n9# in Gnd Gnd nfet w=4 l=2
+  ad=0 pd=0 as=20 ps=18
M1003 out in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in Gnd 0.03fF
C1 vdd in 0.33fF
C2 out Gnd 0.08fF
C3 out vdd 0.58fF
C4 out in 0.11fF
C5 Gnd 0 0.11fF $ **FLOATING
C6 out 0 0.26fF $ **FLOATING
C7 in 0 0.37fF $ **FLOATING
C8 vdd 0 0.55fF $ **FLOATING
