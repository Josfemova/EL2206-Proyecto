magic
tech scmos
timestamp 1667803018
<< nwell >>
rect -17 1 24 26
<< ntransistor >>
rect -6 -9 0 -5
rect 4 -9 10 -5
<< ptransistor >>
rect -3 7 -1 15
rect 5 7 7 15
<< ndiffusion >>
rect -7 -9 -6 -5
rect 0 -9 4 -5
rect 10 -9 11 -5
<< pdiffusion >>
rect -4 7 -3 15
rect -1 7 0 15
rect 4 7 5 15
rect 7 7 8 15
<< ndcontact >>
rect -11 -9 -7 -5
rect 11 -9 15 -5
<< pdcontact >>
rect -8 7 -4 15
rect 0 7 4 15
rect 8 7 12 15
<< psubstratepcontact >>
rect -11 -17 -7 -13
rect 0 -17 4 -13
rect 11 -17 15 -13
<< nsubstratencontact >>
rect -8 19 -4 23
rect 0 19 4 23
rect 8 19 12 23
<< polysilicon >>
rect -3 15 -1 27
rect 5 15 7 27
rect -3 -2 -1 7
rect 5 -2 7 7
rect 18 3 20 27
rect -6 -5 0 -2
rect 4 -5 10 -2
rect -6 -12 0 -9
rect 4 -12 10 -9
rect -3 -19 -1 -12
rect 5 -19 7 -12
rect 18 -19 20 -1
<< polycontact >>
rect -4 27 0 31
rect 4 27 8 31
rect 17 27 21 31
rect 17 -1 21 3
<< metal1 >>
rect -4 31 8 35
rect 17 31 21 35
rect -17 19 -8 23
rect -4 19 0 23
rect 4 19 8 23
rect 12 19 21 23
rect 0 15 4 19
rect -8 3 -4 7
rect 8 3 12 7
rect -11 -1 17 3
rect -11 -5 -7 -1
rect -11 -13 -7 -9
rect -17 -17 -11 -13
rect -7 -17 0 -13
rect 4 -17 11 -13
rect 15 -17 24 -13
<< labels >>
rlabel metal1 0 31 4 35 5 in
rlabel metal1 -14 19 -10 23 3 vdd
rlabel metal1 -15 -17 -11 -13 2 Gnd
rlabel metal1 17 31 21 35 6 out
<< end >>
